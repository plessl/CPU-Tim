module pRom(
    input wire clock,
    input wire ce,
    input wire oce,
    input wire reset,
    addr,
    dataout
);

endmodule